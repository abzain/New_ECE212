//------------------------------------------------
// mipsparts.sv
// David_Harris@hmc.edu 23 October 2005
// Updated to SystemVerilog dmh 12 November 2010
// Components used in MIPS processor
//------------------------------------------------

module regfile(input  logic        clk, 
               input  logic        we3, 
               input  logic [4:0]  ra1, ra2, wa3, 
               input  logic [31:0] wd3, 
               output logic [31:0] rd1, rd2);

  logic [31:0] rf[31:0];

  // three ported register file
  // read two ports combinationally
  // write third port on rising edge of clock
  // register 0 hardwired to 0

  always_ff @(posedge clk)
    if (we3) rf[wa3] <= wd3;	

  assign rd1 = (ra1 != 0) ? rf[ra1] : 0;
  assign rd2 = (ra2 != 0) ? rf[ra2] : 0;
endmodule

module adder(input  logic [31:0] a, b,
             output logic [31:0] y);

  assign y = a + b;
endmodule

module sl2(input  logic [31:0] a,
           output logic [31:0] y);

  // shift left by 2
  assign y = {a[29:0], 2'b00};
endmodule

module signext(input  logic [15:0] a,
               output logic [31:0] y);
              
  assign y = {{16{a[15]}}, a};
endmodule

<<<<<<< HEAD
//ADDED ZERO EXTENDER
module zeroext(input  logic [15:0] a,
               output logic [31:0] y);
              
  assign y = {{16{1'b0}}, a};
=======
//zero extending added
module zeroext(input  logic [15:0] a,
               output logic [31:0] y);
              
  assign y = {16'h0000, a};
>>>>>>> origin/master
endmodule

module flopr #(parameter WIDTH = 8)
              (input  logic             clk, reset,
               input  logic [WIDTH-1:0] d, 
               output logic [WIDTH-1:0] q);

  always_ff @(posedge clk, posedge reset)
    if (reset) q <= 0;
    else       q <= d;
endmodule

module flopenr #(parameter WIDTH = 8)
                (input  logic             clk, reset,
                 input  logic             en,
                 input  logic [WIDTH-1:0] d, 
                 output logic [WIDTH-1:0] q);
 
  always_ff @(posedge clk, posedge reset)
    if      (reset) q <= 0;
    else if (en)    q <= d;
endmodule

module mux2 #(parameter WIDTH = 8)
             (input  logic [WIDTH-1:0] d0, d1, 
              input  logic             s, 
              output logic [WIDTH-1:0] y);
              
   always_comb
     case(s)
         1'b0: y <= d0;
         1'b1: y <= d1;
         default: y <= 8'hxx;
     endcase
endmodule

//MODIFIED MUX TO TAKE EXTRA INPUT              
module mux3 #(parameter WIDTH = 8)
               (input  logic [WIDTH-1:0] d0, d1, k, 
                input  logic [1:0]       s, 
                output logic [WIDTH-1:0] y);

<<<<<<< HEAD
// always_comb
//    case(s)
//        2'b00: y <= d0;
//        2'b01: y <= k;
//        2'b10: y <= d1;
//        default: y <= 6'dx;
//    endcase
=======
     always_comb
        case(s)
            2'b00: y <= d0;
            2'b01: y <= d1;
            2'b10: y <= k;
            default: y <= 8'hxx;
        endcase
>>>>>>> origin/master
endmodule
